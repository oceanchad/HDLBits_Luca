module top_module (
    input clk,
    input reset,            // Synchronous reset
    input [7:0] d,
    output [7:0] q
);
    always_ff@(posedge clk) begin
        if (reset == 1'b1)
            q <= 7'b0;
        else
            q <= d;
    end

endmodule
